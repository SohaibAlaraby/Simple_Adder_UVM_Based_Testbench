interface aintf(input bit clk);// #(parameter bits = 4);
  logic [3 : 0] A;
  logic [3 : 0] B;
  logic [3 : 0] sum;
  logic cout;
    
endinterface:aintf //interfacename
